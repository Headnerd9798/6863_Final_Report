module ALW_NR_TCST (out_a);
   output reg [1:0] out_a;

   always@(posedge 1)
   out_a <= 2'b00;
endmodule
