module VAR_NR_TIME (port_a);
   output port_a;
   time t1;
   assign port_a = t1;
endmodule
