module CST_MS_LPDZ (out_a);
   output [1:0] out_a;
   wire [1:0] wire_a= 1'b0;
   assign out_a = wire_a;
endmodule
