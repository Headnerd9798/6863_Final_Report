module SIG_NR_NDCL (inp, outp);   
   input inp;   
   output outp;
   wor inp;   
   assign outp = inp; 
endmodule

