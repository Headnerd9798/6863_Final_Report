module MOD_NR_FINB (port_a);
   output reg port_a;
   final
   port_a = 1'b0;
endmodule
