module CST_MS_SIZE (outp);
   output outp;
   assign outp = 3'b11111;
endmodule
