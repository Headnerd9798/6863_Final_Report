module MOD_NR_PGAT (a, out1);
   input a;
   output out1;
   buf b1(out1,a);
endmodule
