module OPR_NR_TRNB (port_a);
   output [2:0] port_a;
   wire[2:0] port_a;
   assign port_a = 4'b0011 + 4'b0011;
endmodule
