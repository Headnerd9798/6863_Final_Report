LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY MOD_NO_PRTD IS

END MOD_NO_PRTD;

ARCHITECTURE MOD_NO_PRTD_rtl OF MOD_NO_PRTD IS
    SIGNAL a, b : std_logic;
BEGIN
    a <= b;
END MOD_NO_PRTD_rtl;
