module MOD_NO_PRTD; 
   reg a, b; 
endmodule 
