module IDN_NR_SVKW (port_a, covergroup);
      input port_a;
      output covergroup;

         assign covergroup = port_a;
endmodule
