module VAR_NR_REAL (port_a);
   output port_a;
   real r1;
   assign port_a = r1;
endmodule
