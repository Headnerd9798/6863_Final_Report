module IDN_NR_ESCA (inp_1); 
   input inp_1;
   wire \wir_* ;
   assign \wir_* = inp_1;
endmodule
