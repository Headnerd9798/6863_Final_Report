module WIR_NO_USED (in1, out1);
   input in1;
   output out1;
   reg out1;
   wire g1;
   always @(in1)
   out1 <= in1;
endmodule
