module ALW_NO_EVTS (in_a);
   input in_a;
   reg out_a;
   reg clk;
   always
   begin
      out_a <= in_a;
   end
endmodule
