module VAR_NR_INDL(count);
   output [1:0] count;
   reg [1:0] reg1 = 2'b01;
   assign count = reg1;
endmodule
