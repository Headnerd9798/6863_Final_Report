module IDN_NF_ALCA (port_a, portB);
   input port_a;
   output portB;
   assign portB = port_a;
endmodule
