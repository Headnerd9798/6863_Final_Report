module ASG_NS_TRNB (out1, out2);
   output [7:0] out1;
   output [7:0] out2;
   assign out1 = 9'b110101010;
   assign out2 = 9'b010101010;
endmodule
