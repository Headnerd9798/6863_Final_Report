module ASG_NR_LMSB (out1);
   output [7:0] out1;
   assign out1 = 9'b110101010;
endmodule
