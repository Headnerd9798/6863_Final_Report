library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

ENTITY flags IS
PORT (
dReady                  : OUT std_logic;
dError                  : OUT std_logic;
clk                     : IN std_logic;
set                     : IN std_logic;
reset                   : IN std_logic;
dIn                     : IN std_logic);
END flags;
ARCHITECTURE rtl OF flags IS
SIGNAL dReady_reg             :  std_logic;
SIGNAL dError_reg             :  std_logic;
BEGIN
dReady <= dReady_reg;
dError <= dError_reg;
PROCESS
BEGIN
WAIT UNTIL (clk'EVENT AND clk = '1');
IF (reset = '1') THEN
dReady_reg <= '0';
dError_reg <= '0';
ELSE
IF (set = '1') THEN
dReady_reg <= dIn;
dError_reg <= NOT dIn;
END IF;
END IF;
END PROCESS;
END rtl;


-- -------------------------------------------------------
-- Copyright (c) 2000 Jasper Design Automation, Inc.
--
-- All rights reserved.
--
-- Jasper Design Automation Proprietary and Confidential.
-- -------------------------------------------------------

