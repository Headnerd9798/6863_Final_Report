module MOD_NR_INIB (port_a);
   output reg port_a;
   initial
   port_a = 1'b0;
endmodule
