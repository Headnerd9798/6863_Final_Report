module MOD_IS_RBXE;
   VERI1139 VERI1139();
endmodule
module VERI1139(r, a, y);
   input real r;
   input int a;
   output int y;
endmodule
