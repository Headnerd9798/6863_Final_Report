module CST_NO_BWID (port_a);
   output port_a;
   assign port_a = 'b000000;
endmodule
