module CST_NR_MSBX (in_a, in_b);
   output [3:0] in_a;
   output [7:0] in_b;
   assign in_a = 4'bx1;
   assign in_b = 4'bxx;
endmodule

