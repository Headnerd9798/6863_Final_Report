module WIR_NO_READ (inp_1);
   input inp_1;
   wire wir_a;
   assign wir_a = inp_1;
endmodule
